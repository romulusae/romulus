module lfsr3_28 (/*AUTOARG*/
   // Outputs
   so,
   // Inputs
   si
   ) ;
   output [127:0] so;
   input [127:0]  si;

   wire [7:0] 	  m [15:0];
   wire [7:0] 	  z [15:0];

   assign m[0] = si[7:0];
   assign m[1] = si[15:8];
   assign m[2] = si[23:16];
   assign m[3] = si[31:24];
   assign m[4] = si[39:32];
   assign m[5] = si[47:40];
   assign m[6] = si[55:48];
   assign m[7] = si[63:56];
   assign m[8] = si[71:64];
   assign m[9] = si[79:72];
   assign m[10] = si[87:80];
   assign m[11] = si[95:88];
   assign m[12] = si[103:96];
   assign m[13] = si[111:104];
   assign m[14] = si[119:112];
   assign m[15] = si[127:120];

   assign z[0] =  {m[0] [5:0],m[0] [7] ^ m[0] [5], m[0] [6]^ m[0][4]};
   assign z[1] =  {m[1] [5:0],m[1] [7] ^ m[1] [5], m[1] [6]^ m[1][4]};
   assign z[2] =  {m[2] [5:0],m[2] [7] ^ m[2] [5], m[2] [6]^ m[2][4]};
   assign z[3] =  {m[3] [5:0],m[3] [7] ^ m[3] [5], m[3] [6]^ m[3][4]};
   assign z[4] =  {m[4] [5:0],m[4] [7] ^ m[4] [5], m[4] [6]^ m[4][4]};
   assign z[5] =  {m[5] [5:0],m[5] [7] ^ m[5] [5], m[5] [6]^ m[5][4]};
   assign z[6] =  {m[6] [5:0],m[6] [7] ^ m[6] [5], m[6] [6]^ m[6][4]};
   assign z[7] =  {m[7] [5:0],m[7] [7] ^ m[7] [5], m[7] [6]^ m[7][4]};
   assign z[8] =  {m[8] [5:0],m[8] [7] ^ m[8] [5], m[8] [6]^ m[8][4]};
   assign z[9] =  {m[9] [5:0],m[9] [7] ^ m[9] [5], m[9] [6]^ m[9][4]};
   assign z[10] = {m[10][5:0],m[10][7] ^ m[10][5], m[10][6]^ m[10][4]};
   assign z[11] = {m[11][5:0],m[11][7] ^ m[11][5], m[11][6]^ m[11][4]};
   assign z[12] = {m[12][5:0],m[12][7] ^ m[12][5], m[12][6]^ m[12][4]};
   assign z[13] = {m[13][5:0],m[13][7] ^ m[13][5], m[13][6]^ m[13][4]};
   assign z[14] = {m[14][5:0],m[14][7] ^ m[14][5], m[14][6]^ m[14][4]};
   assign z[15] = {m[15][5:0],m[15][7] ^ m[15][5], m[15][6]^ m[15][4]};

   assign so = {z[15],
		z[14],
		z[13],
		z[12],
		z[11],
		z[10],
		z[9],
		z[8],
		z[7],
		z[6],
		z[5],
		z[4],
		z[3],
		z[2],
		z[1],
		z[0]};
   
   
   
   
endmodule // lfsr2_38
